    `define PRESCALE_W      24
    `define ADDR_W          5
    `define DATA_W          10