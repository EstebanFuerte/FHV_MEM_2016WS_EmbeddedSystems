// ------------------------------------
// MEM3 -- HDL
// Project:		
// Author:		stst
// Date:		30.01.2017
// ------------------------------------

module sevenseg(
	// Define inputs and outputs
);

	always_comb begin
		
	end
	
	// outside an always - assign is necessary
	

endmodule